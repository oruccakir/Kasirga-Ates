// Purpose: Control Unit for the Execute stage of the pipeline.
// Functionality: This module performs the control of the pipeline.
// File: ControlUnit.v

module ControlUnit (
    input wire clk_i, // Clock input
    input wire rst_i, // Reset input
);


endmodule
