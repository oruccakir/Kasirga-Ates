// Purpose: Memory step module for the pipeline.
// Functionality: This module performs the memory stage of the pipeline.
// File: MemoryStep.v

module MemoryStep (
    input wire clk_i, // Clock input
    input wire rst_i, // Reset input
);
    

endmodule