// Purpose: Execute Step 1 of the pipeline.
// Functionality: This module performs the first part of the execute stage of the pipeline.
// File: ExecuteStep1.v

module ExecuteStep1 (
    input wire clk_i, // Clock input
    input wire rst_i, // Reset input
);
    

endmodule