// Purpose: Processor module for the pipeline processor.
// Functional Description: This module is the main module for the processor. It is responsible for the execution of the instructions. It is also responsible for the control signals of the pipeline.
// File: Processor.v

// Include the definitions
`include "definitions.v"

module Processor(
    input wire clk_i,
    input wire rst_i,
    input wire [31:0] mem_address_i,
);

endmodule
