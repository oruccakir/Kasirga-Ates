// File: definitions.vh
// Purpose: Contains definitions for the pipeline processor.

// CONTROL SIGNALS FOR REGISTER FILE SELECTION
`define INTEGER_REGISTER        2'b0
`define FLOAT_REGISTER          2'b1
`define CSR_REGISTER            2'b10

// CONTROL SIGNALS FOR UNIT SELECTION 
`define FLOATING_POINT_UNIT             4'h0
`define ARITHMETIC_LOGIC_UNIT           4'h1
`define INTEGER_MULTIPLICATION_UNIT     4'h2
`define INTEGER_DIVISION_UNIT           4'h3
`define BRANCH_RESOLVER_UNIT            4'h4
`define CONTROL_UNIT                    4'h5
`define CONTROL_STATUS_UNIT             4'h6
`define ATOMIC_UNIT                     4'h7
`define BIT_MANIPULATION_UNIT           4'h8
`define MEMORY_UNIT                     4'h9


// Control Signals for ALU operations
`define ALU_ADD                 5'h0
`define ALU_SUB                 5'h1
`define ALU_XOR                 5'h2
`define ALU_OR                  5'h3
`define ALU_AND                 5'h4
`define ALU_SLL                 5'h5
`define ALU_SRL                 5'h6
`define ALU_SRA                 5'h7
`define ALU_SLT                 5'h8
`define ALU_SLTU                5'h9
`define ALU_ADDI                5'ha
`define ALU_SLTI                5'hb
`define ALU_SLTIU               5'hc
`define ALU_XORI                5'hd
`define ALU_ORI                 5'he
`define ALU_ANDI                5'hf
`define ALU_SLLI                5'h10
`define ALU_SRLI                5'h11
`define ALU_SRAI                5'h12
`define ALU_SRLI                5'h13
`define ALU_SRAI                5'h14
`define ALU_AUIPC               5'h15
`define ALU_LUI                 5'h16

// Control Signals integer multiplication and division operations
`define INT_MUL                 4'h0
`define INT_MULH                4'h1
`define INT_MULHSU              4'h2
`define INT_MULHU               4'h3
`define INT_DIV                 4'h4
`define INT_DIVU                4'h5
`define INT_REM                 4'h6
`define INT_REMU                4'h7


// Control Signals for Atomic operations
`define ATOM_LR_W               4'h0
`define ATOM_SC_W               4'h1
`define ATOM_AMOSWAP_W          4'h2
`define ATOM_AMOADD_W           4'h3
`define ATOM_AMOXOR_W           4'h4
`define ATOM_AMOAND_W           4'h5
`define ATOM_AMOOR_W            4'h6
`define ATOM_AMOMIN_W           4'h7
`define ATOM_AMOMAX_W           4'h8
`define ATOM_AMOMINU_W          4'h9
`define ATOM_AMOMAXU_W          4'hA

// Control Signals for floating point operations
`define FLT_FLW                5'h0
`define FLT_FSW                5'h1
`define FLT_FMADD_S            5'h2
`define FLT_FMSUB_S            5'h3
`define FLT_FNMSUB_S           5'h4
`define FLT_FNMADD_S           5'h5
`define FLT_FADD_S             5'h6
`define FLT_FSUB_S             5'h7
`define FLT_FMUL_S             5'h8
`define FLT_FDIV_S             5'h9
`define FLT_FSQRT_S            5'hA
`define FLT_FSGNJ_S            5'hB
`define FLT_FSGNJN_S           5'hC
`define FLT_FSGNJX_S           5'hD
`define FLT_FMIN_S             5'hE
`define FLT_FMAX_S             5'hF
`define FLT_FCVT_W_S           5'h10
`define FLT_FCVT_WU_S          5'h11
`define FLT_FMV_X_W            5'h12
`define FLT_FEQ_S              5'h13
`define FLT_FLT_S              5'h14
`define FLT_FLE_S              5'h15
`define FLT_FCLASS_S           5'h16
`define FLT_FCVT_S_W           5'h17
`define FLT_FCVT_S_WU          5'h18
`define FLT_FMV_W_X            5'h19

// Control Signals for bit manipulation operations
`define BT_ANDN                 5'h0
`define BT_CLMUL                5'h1
`define BT_CLMULH               5'h2
`define BT_CLMULR               5'h3
`define BT_CLZ                  5'h4
`define BT_CPOP                 5'h5
`define BT_CTZ                  5'h6
`define BT_MAX                  5'h7
`define BT_MAXU                 5'h8
`define BT_MIN                  5'h9
`define BT_MINU                 5'hA
`define BT_ORC_B                5'hB
`define BT_ORN                  5'hC
`define BT_REV8                 5'hD
`define BT_ROL                  5'hE
`define BT_ROR                  5'hF
`define BT_RORI                 5'h10
`define BT_BCLR                 5'h11
`define BT_BCLRI                5'h12
`define BT_BEXT                 5'h13
`define BT_BEXTI                5'h14
`define BT_BINV                 5'h15
`define BT_BINVI                5'h16
`define BT_BSET                 5'h17
`define BT_BSETI                5'h18
`define BT_SEXT_B               5'h19
`define BT_SEXT_H               5'h1A
`define BT_SH1ADD               5'h1B
`define BT_SH2ADD               5'h1C
`define BT_SH3ADD               5'h1D
`define BT_XNOR                 5'h1E
`define BT_ZEXT_H               5'h1F


// For memory instructions
`define MEM_LB                          3'h0
`define MEM_LH                          3'h1
`define MEM_LW                          3'h2
`define MEM_LBU                         3'h3
`define MEM_LHU                         3'h4
`define MEM_SB                          3'h5
`define MEM_SH                          3'h6
`define MEM_SW                          3'h7

// Control Signals For Branch Resolver Unit
`define BR_BEQ                          3'h0
`define BR_BNE                          3'h1
`define BR_BLT                          3'h2
`define BR_BGE                          3'h3
`define BR_BLTU                         3'h4
`define BR_BGEU                         3'h5
`define BR_JAL                          3'h6
`define BR_JALR                         3'h7


// Control Signals for Memory operations //sebebi bilinmiyor
// for integer memory operations
`define MEM_LOAD                3'b000
`define MEM_STORE               3'b001
// for floating point memory operations
`define FMEM_LOAD               3'b010
`define FMEM_STORE              3'b011
// for atomic memory operations
`define ATOM_MEM_LOAD           3'b100
`define ATOM_MEM_STORE          3'b101

//RV32I Buyruklari
`define ADD         32'b0000000_?????_?????_000_?????_0110011
`define SUB         32'b0100000_?????_?????_000_?????_0110011
`define SLL         32'b0000000_?????_?????_001_?????_0110011
`define SLT         32'b0000000_?????_?????_010_?????_0110011
`define SLTU        32'b0000000_?????_?????_011_?????_0110011
`define XOR         32'b0000000_?????_?????_100_?????_0110011
`define SRL         32'b0000000_?????_?????_101_?????_0110011
`define SRA         32'b0100000_?????_?????_101_?????_0110011
`define OR          32'b0000000_?????_?????_110_?????_0110011
`define AND         32'b0000000_?????_?????_111_?????_0110011

`define ADDI        32'b????????????_?????_000_?????_0010011
`define SLTI        32'b????????????_?????_010_?????_0010011
`define SLTIU       32'b????????????_?????_011_?????_0010011
`define XORI        32'b????????????_?????_100_?????_0010011
`define ORI         32'b????????????_?????_110_?????_0010011
`define ANDI        32'b????????????_?????_111_?????_0010011

`define SLLI        32'b0000000_?????_?????_001_?????_0010011
`define SRLI        32'b0000000_?????_?????_101_?????_0010011
`define SRAI        32'b0100000_?????_?????_101_?????_0010011

`define SB          32'b???????_?????_?????_000_?????_0100011
`define SH          32'b???????_?????_?????_001_?????_0100011
`define SW          32'b???????_?????_?????_010_?????_0100011

`define LB          32'b????????????_?????_000_?????_0000011
`define LH          32'b????????????_?????_001_?????_0000011
`define LW          32'b????????????_?????_010_?????_0000011
`define LBU         32'b????????????_?????_100_?????_0000011
`define LHU         32'b????????????_?????_101_?????_0000011

`define BEQ         32'b?_??????_?????_?????_000_????_?_1100011
`define BNE         32'b?_??????_?????_?????_001_????_?_1100011
`define BLT         32'b?_??????_?????_?????_100_????_?_1100011
`define BGE         32'b?_??????_?????_?????_101_????_?_1100011
`define BLTU        32'b?_??????_?????_?????_110_????_?_1100011
`define BGEU        32'b?_??????_?????_?????_111_????_?_1100011

`define LUI         32'b????????????????????_?????_0110111
`define AUIPC       32'b????????????????????_?????_0010111

`define JAL         32'b?_??????????_?_????????_?????_0010111
`define JALR        32'b?_??????????_?_????????_?????_0010111

//RV32M Buyruklari
`define MUL         32'b0000001_?????_?????_000_?????_0110011
`define MULH        32'b0000001_?????_?????_001_?????_0110011
`define MULHSU      32'b0000001_?????_?????_010_?????_0110011
`define MULHU       32'b0000001_?????_?????_011_?????_0110011
`define DIV         32'b0000001_?????_?????_100_?????_0110011
`define DIVU        32'b0000001_?????_?????_101_?????_0110011
`define REM         32'b0000001_?????_?????_110_?????_0110011
`define REMU        32'b0000001_?????_?????_111_?????_0110011


//RV32A Buyruklari
`define LR_W        32'b00010_?_?_00000_?????_010_?????_0101111
`define SC_W        32'b00011_?_?_?????_?????_010_?????_0101111
`define AMOSWAP_W   32'b00001_?_?_?????_?????_010_?????_0101111
`define AMOADD_W    32'b00000_?_?_?????_?????_010_?????_0101111
`define AMOXOR_W    32'b00100_?_?_?????_?????_010_?????_0101111
`define AMOAND_W    32'b01100_?_?_?????_?????_010_?????_0101111
`define AMOOR_W     32'b01000_?_?_?????_?????_010_?????_0101111
`define AMOMIN_W    32'b10000_?_?_?????_?????_010_?????_0101111
`define AMOMAX_W    32'b10100_?_?_?????_?????_010_?????_0101111
`define AMOMINU_W   32'b11000_?_?_?????_?????_010_?????_0101111
`define AMOMAXU_W   32'b11100_?_?_?????_?????_010_?????_0101111

//RV32F Buyruklari
`define FLW         32'b????????????_?????_010_?????_0000111
`define FSW         32'b???????_?????_?????_010_?????_0100111
`define FMADD_S     32'b?????_00_?????_?????_???_?????_1000011
`define FMSUB_S     32'b?????_00_?????_?????_???_?????_1000111
`define FNMSUB_S    32'b?????_00_?????_?????_???_?????_1001011
`define FNMADD_S    32'b?????_00_?????_?????_???_?????_1001111
`define FADD_S      32'b0000000_?????_?????_???_?????_1010011
`define FSUB_S      32'b0000100_?????_?????_???_?????_1010011
`define FMUL_S      32'b0001000_?????_?????_???_?????_1010011
`define FDIV_S      32'b0101100_?????_?????_???_?????_1010011
`define FSQRT_S     32'b0101100_00000_?????_???_?????_1010011
`define FSGNJ_S     32'b0010000_?????_?????_000_?????_1010011
`define FSGNJN_S    32'b0010000_?????_?????_001_?????_1010011
`define FSGNJX_S    32'b0010000_?????_?????_010_?????_1010011
`define FMIN_S      32'b0010100_?????_?????_000_?????_1010011
`define FMAX_S      32'b0010100_?????_?????_001_?????_1010011
`define FCVT_W_S    32'b1100000_00000_?????_???_?????_1010011
`define FCVT_WU_S   32'b1100000_00001_?????_???_?????_1010011
`define FMV_X_W     32'b1110000_00000_?????_000_?????_1010011
`define FEQ_S       32'b1010000_?????_?????_010_?????_1010011
`define FLT_S       32'b1010000_?????_?????_001_?????_1010011
`define FLE_S       32'b1010000_?????_?????_000_?????_1010011
`define FCLASS_S    32'b1110000_00000_?????_001_?????_1010011
`define FCVT_S_W    32'b1101000_00000_?????_???_?????_1010011
`define FCVT_S_WU   32'b1101000_00001_?????_???_?????_1010011
`define FMV_W_X     32'b1111000_00000_?????_000_?????_1010011

//RV32B Buyruklari
`define ANDN        32'b0100000_?????_?????_111_?????_0110011
`define CLMUL       32'b0000101_?????_?????_001_?????_0110011
`define CLMULH      32'b0000101_?????_?????_011_?????_0110011
`define CLMULR      32'b0000101_?????_?????_010_?????_0110011
`define CLZ         32'b0110000_00000_?????_001_?????_0010011
`define CPOP        32'b0110000_00010_?????_001_?????_0010011
`define CTZ         32'b0110000_00010_?????_001_?????_0010011
`define MAX         32'b0000101_?????_?????_110_?????_0110011
`define MAXU        32'b0000101_?????_?????_111_?????_0110011
`define MIN         32'b0000101_?????_?????_100_?????_0110011
`define MINU        32'b0000101_?????_?????_101_?????_0110011
`define ORC_B       32'b0010100_00111_?????_101_?????_0010011
`define ORN         32'b0100000_?????_?????_110_?????_0110011
`define REV8        32'b0110100_11000_?????_101_?????_0010011
`define ROL         32'b0110000_?????_?????_001_?????_0110011
`define ROR         32'b0110000_?????_?????_101_?????_0110011
`define RORI        32'b0110000_?????_?????_101_?????_0010011
`define BCLR        32'b0100100_?????_?????_001_?????_0110011
`define BCLRI       32'b0100100_?????_?????_001_?????_0010011
`define BEXT        32'b0100100_?????_?????_101_?????_0110011
`define BEXTI       32'b0100100_?????_?????_101_?????_0010011
`define BINV        32'b0110100_?????_?????_001_?????_0110011
`define BINVI       32'b0110100_?????_?????_001_?????_0010011
`define BSET        32'b0010100_?????_?????_001_?????_0110011
`define BSETI       32'b0010100_?????_?????_001_?????_0010011
`define SEXT_B      32'b0110000_00100_?????_001_?????_0010011
`define SEXT_H      32'b0110000_00101_?????_001_?????_0010011
`define SH1ADD      32'b0010000_?????_?????_010_?????_0110011
`define SH2ADD      32'b0010000_?????_?????_100_?????_0110011
`define SH3ADD      32'b0010000_?????_?????_110_?????_0110011
`define XNOR        32'b0100000_?????_?????_100_?????_0110011
`define ZEXT_H      32'b0000100_00000_?????_100_?????_0110011


// Buyrukların çözülmesi için gereken bitler(Bit manipülasyon buyrukları eklenerek en düşük bit sayısı ve değerli bitler bulunarak oluşturulacaktır) 
`define BIT_SAYISI_COZ 19 //(31-27, 25-20, 14-12, 6-2)

`define ADD_COZ            19'b000000?????00001100
`define SUB_COZ            19'b010000?????00001100
`define SLL_COZ            19'b000000?????00101100
`define SLT_COZ            19'b000000?????01001100
`define SLTU_COZ           19'b000000?????01101100
`define XOR_COZ            19'b000000?????10001100
`define SRL_COZ            19'b000000?????10101100
`define SRA_COZ            19'b010000?????10101100
`define OR_COZ             19'b000000?????11001100
`define AND_COZ            19'b000000?????11101100
`define ADDI_COZ           19'b???????????00000100
`define SLTI_COZ           19'b???????????01000100
`define SLTIU_COZ          19'b???????????01100100
`define XORI_COZ           19'b???????????10000100
`define ORI_COZ            19'b???????????11000100
`define ANDI_COZ           19'b???????????11100100
`define SLLI_COZ           19'b000000?????00100100
`define SRLI_COZ           19'b000000?????10100100
`define SRAI_COZ           19'b010000?????10100100
`define SB_COZ             19'b???????????00001000
`define SH_COZ             19'b???????????00101000
`define SW_COZ             19'b???????????01001000
`define LB_COZ             19'b???????????00000000
`define LH_COZ             19'b???????????00100000
`define LW_COZ             19'b???????????01000000
`define LBU_COZ            19'b???????????10000000
`define LHU_COZ            19'b???????????10100000
`define BEQ_COZ            19'b???????????00011000
`define BNE_COZ            19'b???????????00111000
`define BLT_COZ            19'b???????????10011000
`define BGE_COZ            19'b???????????10111000
`define BLTU_COZ           19'b???????????11011000
`define BGEU_COZ           19'b???????????11111000
`define LUI_COZ            19'b??????????????01101
`define AUIPC_COZ          19'b??????????????00101
`define JAL_COZ            19'b??????????????00101
`define JALR_COZ           19'b??????????????00101
`define MUL_COZ            19'b000001?????00001100
`define MULH_COZ           19'b000001?????00101100
`define MULHSU_COZ         19'b000001?????01001100
`define MULHU_COZ          19'b000001?????01101100
`define DIV_COZ            19'b000001?????10001100
`define DIVU_COZ           19'b000001?????10101100
`define REM_COZ            19'b000001?????11001100
`define REMU_COZ           19'b000001?????11101100
`define LR_W_COZ           19'b00010?0000001001011
`define SC_W_COZ           19'b00011??????01001011
`define AMOSWAP_W_COZ      19'b00001??????01001011
`define AMOADD_W_COZ       19'b00000??????01001011
`define AMOXOR_W_COZ       19'b00100??????01001011
`define AMOAND_W_COZ       19'b01100??????01001011
`define AMOOR_W_COZ        19'b01000??????01001011
`define AMOMIN_W_COZ       19'b10000??????01001011
`define AMOMAX_W_COZ       19'b10100??????01001011
`define AMOMINU_W_COZ      19'b11000??????01001011
`define AMOMAXU_W_COZ      19'b11100??????01001011
`define FLW_COZ            19'b???????????01000001
`define FSW_COZ            19'b???????????01001001
`define FMADD_S_COZ        19'b?????0????????10000
`define FMSUB_S_COZ        19'b?????0????????10001
`define FNMSUB_S_COZ       19'b?????0????????10010
`define FNMADD_S_COZ       19'b?????0????????10011
`define FADD_S_COZ         19'b000000????????10100
`define FSUB_S_COZ         19'b000010????????10100
`define FMUL_S_COZ         19'b000100????????10100
`define FDIV_S_COZ         19'b010110????????10100
`define FSQRT_S_COZ        19'b01011000000???10100
`define FSGNJ_S_COZ        19'b001000?????00010100
`define FSGNJN_S_COZ       19'b001000?????00110100
`define FSGNJX_S_COZ       19'b001000?????01010100
`define FMIN_S_COZ         19'b001010?????00010100
`define FMAX_S_COZ         19'b001010?????00110100
`define FCVT_W_S_COZ       19'b11000000000???10100
`define FCVT_WU_S_COZ      19'b11000000001???10100
`define FMV_X_W_COZ        19'b1110000000000010100
`define FEQ_S_COZ          19'b101000?????01010100
`define FLT_S_COZ          19'b101000?????00110100
`define FLE_S_COZ          19'b101000?????00010100
`define FCLASS_S_COZ       19'b1110000000000110100
`define FCVT_S_W_COZ       19'b11010000000???10100
`define FCVT_S_WU_COZ      19'b11010000001???10100
`define FMV_W_X_COZ        19'b1111000000000010100
`define ANDN_COZ           19'b010000?????11101100
`define CLMUL_COZ          19'b000011?????00101100
`define CLMULH_COZ         19'b000011?????01101100
`define CLMULR_COZ         19'b000011?????01001100
`define CLZ_COZ            19'b0110000000000100100
`define CPOP_COZ           19'b0110000001000100100
`define CTZ_COZ            19'b0110000001000100100
`define MAX_COZ            19'b000011?????11001100
`define MAXU_COZ           19'b000011?????11101100
`define MIN_COZ            19'b000011?????10001100
`define MINU_COZ           19'b000011?????10101100
`define ORC_B_COZ          19'b0010100011110100100
`define ORN_COZ            19'b010000?????11001100
`define REV8_COZ           19'b0110101100010100100
`define ROL_COZ            19'b011000?????00101100
`define ROR_COZ            19'b011000?????10101100
`define RORI_COZ           19'b011000?????10100100
`define BCLR_COZ           19'b010010?????00101100
`define BCLRI_COZ          19'b010010?????00100100
`define BEXT_COZ           19'b010010?????10101100
`define BEXTI_COZ          19'b010010?????10100100
`define BINV_COZ           19'b011010?????00101100
`define BINVI_COZ          19'b011010?????00100100
`define BSET_COZ           19'b001010?????00101100
`define BSETI_COZ          19'b001010?????00100100
`define SEXT_B_COZ         19'b0110000010000100100
`define SEXT_H_COZ         19'b0110000010100100100
`define SH1ADD_COZ         19'b001000?????01001100
`define SH2ADD_COZ         19'b001000?????10001100
`define SH3ADD_COZ         19'b001000?????11001100
`define XNOR_COZ           19'b010000?????10001100
`define ZEXT_H_COZ         19'b0000100000010001100 



