// Purpose: WriteBackStep module for the WriteBack stage of the pipeline.
// Functionality: This module performs the write back stage of the pipeline.
// File: WriteBackStep.v

module WriteBackStep (
    input wire clk_i, // Clock input
    input wire rst_i, // Reset input
);
    

endmodule