// File: definitions.vh
// Purpose: Contains definitions for the pipeline processor.

// Control Signals for ALU operations
`define ALU_ADDITION = 4'h0
`define ALU_SUBTRACTION = 4'h1
`define ALU_XOR = 4'h2
`define ALU_OR = 4'h3
`define ALU_AND = 4'h4
`define ALU_SLL = 4'h5
`define ALU_SRL = 4'h6
`define ALU_SRA = 4'h7
`define ALU_SLT = 4'h8
`define ALU_SLTU = 4'h9